Holmes Rangemaster Plots

.lib ../../germaniumbjts.lib holmes2017

.include rangemaster.mod

.param vol=0.99

X1 in out rangemaster vol=vol

.param amp=1
.param frq=440

Vin in 0 sin(0 {amp} {frq} 0 0)

.control
foreach ampi 0.1 0.5 1
  alterparam amp=$ampi
  foreach frqi 200
    alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 200Hz input signal
tran 22.675u 0.12 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-rangemaster v(out)

  end
  foreach frqi 500
    alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 500Hz input signal
tran 22.675u 0.108 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-rangemaster v(out)

  end
  foreach frqi 1200
    alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 1200Hz input signal
tran 22.675u 0.103 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-rangemaster v(out)

  end
end
.endc

.end
