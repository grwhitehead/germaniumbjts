Holmes Fuzz Face Plots

.lib ../../germaniumbjts.lib holmes2017

.include fuzzface.mod

.param fuz=0.99
.param vol=0.99

X1 in out fuzzface fuz=fuz vol=vol

.param amp=1
.param frq=440

Vin in 0 sin(0 {amp} {frq} 0 0)

.control
foreach fuzi 0.01 0.1 0.5 0.99
  alterparam fuz=$fuzi
  foreach ampi 0.001 0.01 0.1
    alterparam amp=$ampi
    foreach frqi 200
      alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 200Hz input signal
tran 22.675u 0.12 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-fuzzface-fuz_{$fuzi} v(out)

    end
    foreach frqi 500
      alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 500Hz input signal
tran 22.675u 0.108 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-fuzzface-fuz_{$fuzi} v(out)

    end
    foreach frqi 1200
      alterparam frq=$frqi

reset
* 44100Hz sampling frequency, capture 4 cycles of 1200Hz input signal
tran 22.675u 0.103 0.100
wrdata data/sin_{$frqi}-amp_{$ampi}-fuzzface-fuz_{$fuzi} v(out)

    end
  end
end
.endc

.end
