Holmes AC128 Plots

.lib ../../germaniumbjts.lib holmes2017

Q1 2 1 0 AC128

.param ib=0

Ib 1 0 DC {ib}
Vce 2 0 DC 0

.control

* Replicate Holmes plot
foreach ibi 75u 501u 750u 1000u
alterparam ib=$ibi
reset
dc Vce -5 5 0.1
wrdata output-ib_{$ibi} i(Vce)
end

* Replicate datasheet plot
dc Vce -5 5 0.1 Ib 1m 10m 1m
wrdata output2 i(Vce)

.endc

.end
